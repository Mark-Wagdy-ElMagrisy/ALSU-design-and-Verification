package enum_pkg;
typedef enum {OR, XOR, ADD, MULT, SHIFT, ROTATE, INVALID_6, INVALID_7} my_opcode;
endpackage
